-- Maheen Shoaib & Jessica Persaud
-- ECE 124
-- Section 201

library ieee;
use ieee.std_logic_1164.all;

-- This code defines a multiplexer that selects one of four 4-bit inputs based on a 2-bit select signal.

entity hex_mux is
port (
    hex_num3, hex_num2, hex_num1, hex_num0 : in std_logic_vector(3 downto 0);  -- Four 4-bit inputs
    mux_select                            : in std_logic_vector(1 downto 0);  -- 2-bit multiplexer select signal
    hex_out                               : out std_logic_vector(3 downto 0)  -- 4-bit multiplexer output
);

end hex_mux;

architecture mux_logic of hex_mux is

begin
    -- Multiplexing logic based on mux_select value
    with mux_select(1 downto 0) select
        hex_out <= hex_num0 when "00",  -- Select hex_num0 when select is "00"
                   hex_num1 when "01",  -- Select hex_num1 when select is "01"
                   hex_num2 when "10",  -- Select hex_num2 when select is "10"
                   hex_num3 when "11";  -- Select hex_num3 when select is "11"
                    
end mux_logic;